
`timescale 1 ns / 1 ps


	module myip_v1_0 #
	(
		// Users to add parameters here
		//(lab10) Users to add parameters here
		parameter CNT_BIT = 31,
		//(lab12)
		parameter integer MEM_IN_0_DATA_WIDTH = 32,
		parameter integer MEM_IN_0_ADDR_WIDTH = 9,
		parameter integer MEM_IN_1_DATA_WIDTH = 32,
		parameter integer MEM_IN_1_ADDR_WIDTH = 9,
		parameter integer MEM_IN_2_DATA_WIDTH = 32,
		parameter integer MEM_IN_2_ADDR_WIDTH = 9,
		parameter integer MEM_IN_3_DATA_WIDTH = 32,
		parameter integer MEM_IN_3_ADDR_WIDTH = 9,
		parameter integer MEM_IN_4_DATA_WIDTH = 32,
		parameter integer MEM_IN_4_ADDR_WIDTH = 9,
		parameter integer MEM_IN_5_DATA_WIDTH = 32,
		parameter integer MEM_IN_5_ADDR_WIDTH = 9,
		parameter integer MEM_IN_6_DATA_WIDTH = 32,
		parameter integer MEM_IN_6_ADDR_WIDTH = 9,
		parameter integer MEM_IN_7_DATA_WIDTH = 32,
		parameter integer MEM_IN_7_ADDR_WIDTH = 9,
		parameter integer MEM_IN_8_DATA_WIDTH = 32,
		parameter integer MEM_IN_8_ADDR_WIDTH = 9,
		parameter integer MEM_IN_9_DATA_WIDTH = 32,
		parameter integer MEM_IN_9_ADDR_WIDTH = 9,
		parameter integer MEM_IN_10_DATA_WIDTH = 32,
		parameter integer MEM_IN_10_ADDR_WIDTH = 9,
		parameter integer MEM_IN_11_DATA_WIDTH = 32,
		parameter integer MEM_IN_11_ADDR_WIDTH = 9,
		parameter integer MEM_IN_12_DATA_WIDTH = 32,
		parameter integer MEM_IN_12_ADDR_WIDTH = 9,
		parameter integer MEM_IN_13_DATA_WIDTH = 32,
		parameter integer MEM_IN_13_ADDR_WIDTH = 9,
		parameter integer MEM_IN_14_DATA_WIDTH = 32,
		parameter integer MEM_IN_14_ADDR_WIDTH = 9,
		parameter integer MEM_IN_15_DATA_WIDTH = 32,
		parameter integer MEM_IN_15_ADDR_WIDTH = 9,
		parameter integer MEM_OUT_0_DATA_WIDTH = 32,
		parameter integer MEM_OUT_0_ADDR_WIDTH = 9,
		parameter integer MEM_OUT_1_DATA_WIDTH = 32,
		parameter integer MEM_OUT_1_ADDR_WIDTH = 9,
		parameter integer MEM_OUT_2_DATA_WIDTH = 32,
		parameter integer MEM_OUT_2_ADDR_WIDTH = 9,
		parameter integer MEM_OUT_3_DATA_WIDTH = 32,
		parameter integer MEM_OUT_3_ADDR_WIDTH = 9,
		parameter integer MEM_OUT_4_DATA_WIDTH = 32,
		parameter integer MEM_OUT_4_ADDR_WIDTH = 9,
		parameter integer MEM_OUT_5_DATA_WIDTH = 32,
		parameter integer MEM_OUT_5_ADDR_WIDTH = 9,
		parameter integer MEM_OUT_6_DATA_WIDTH = 32,
		parameter integer MEM_OUT_6_ADDR_WIDTH = 9,
		parameter integer MEM_OUT_7_DATA_WIDTH = 32,
		parameter integer MEM_OUT_7_ADDR_WIDTH = 9,
		parameter integer MEM_OUT_8_DATA_WIDTH = 32,
		parameter integer MEM_OUT_8_ADDR_WIDTH = 9,
		parameter integer MEM_OUT_9_DATA_WIDTH = 32,
		parameter integer MEM_OUT_9_ADDR_WIDTH = 9,
		parameter integer MEM_OUT_10_DATA_WIDTH = 32,
		parameter integer MEM_OUT_10_ADDR_WIDTH = 9,
		parameter integer MEM_OUT_11_DATA_WIDTH = 32,
		parameter integer MEM_OUT_11_ADDR_WIDTH = 9,
		parameter integer MEM_OUT_12_DATA_WIDTH = 32,
		parameter integer MEM_OUT_12_ADDR_WIDTH = 9,
		parameter integer MEM_OUT_13_DATA_WIDTH = 32,
		parameter integer MEM_OUT_13_ADDR_WIDTH = 9,
		parameter integer MEM_OUT_14_DATA_WIDTH = 32,
		parameter integer MEM_OUT_14_ADDR_WIDTH = 9,
		parameter integer MEM_OUT_15_DATA_WIDTH = 32,
		parameter integer MEM_OUT_15_ADDR_WIDTH = 9,
		parameter integer MEM_OUT_16_DATA_WIDTH = 32,
		parameter integer MEM_OUT_16_ADDR_WIDTH = 9,
		parameter integer MEM_OUT_17_DATA_WIDTH = 32,
		parameter integer MEM_OUT_17_ADDR_WIDTH = 9,

		// User parameters ends
		// Do not modify the parameters beyond this line
		// Parameters of Axi Slave Bus Interface S00_AXI
		parameter integer C_S00_AXI_DATA_WIDTH	= 32,
		parameter integer C_S00_AXI_ADDR_WIDTH	= 9
	)
	(
		// Memory I/F
		// Input Bram	
		output		[MEM_IN_0_ADDR_WIDTH-1:0] 	mem_in_0_addr1,
		output		 							mem_in_0_ce1,
		output		 							mem_in_0_we1,
		input 		[MEM_IN_0_DATA_WIDTH-1:0] 	mem_in_0_q1,
		output		[MEM_IN_0_DATA_WIDTH-1:0] 	mem_in_0_d1,
		
		output		[MEM_IN_1_ADDR_WIDTH-1:0] 	mem_in_1_addr1,
		output		 							mem_in_1_ce1,
		output		 							mem_in_1_we1,
		input 		[MEM_IN_1_DATA_WIDTH-1:0]	mem_in_1_q1,
		output		[MEM_IN_1_DATA_WIDTH-1:0] 	mem_in_1_d1,
		
		output		[MEM_IN_2_ADDR_WIDTH-1:0] 	mem_in_2_addr1,
		output		 							mem_in_2_ce1,
		output		 							mem_in_2_we1,
		input 		[MEM_IN_2_DATA_WIDTH-1:0] 	mem_in_2_q1,
		output		[MEM_IN_2_DATA_WIDTH-1:0] 	mem_in_2_d1,
		
		output		[MEM_IN_3_ADDR_WIDTH-1:0] 	mem_in_3_addr1,
		output		 							mem_in_3_ce1,
		output		 							mem_in_3_we1,
		input 		[MEM_IN_3_DATA_WIDTH-1:0]   mem_in_3_q1,
		output		[MEM_IN_3_DATA_WIDTH-1:0] 	mem_in_3_d1,
		
		output		[MEM_IN_4_ADDR_WIDTH-1:0] 	mem_in_4_addr1,
		output		 							mem_in_4_ce1,
		output		 							mem_in_4_we1,
		input 		[MEM_IN_4_DATA_WIDTH-1:0]   mem_in_4_q1,
		output		[MEM_IN_4_DATA_WIDTH-1:0] 	mem_in_4_d1,
		
		output		[MEM_IN_5_ADDR_WIDTH-1:0] 	mem_in_5_addr1,
		output		 							mem_in_5_ce1,
		output		 							mem_in_5_we1,
		input 		[MEM_IN_5_DATA_WIDTH-1:0]   mem_in_5_q1,
		output		[MEM_IN_5_DATA_WIDTH-1:0] 	mem_in_5_d1,
		
		output		[MEM_IN_6_ADDR_WIDTH-1:0] 	mem_in_6_addr1,
		output		 							mem_in_6_ce1,
		output		 							mem_in_6_we1,
		input 		[MEM_IN_6_DATA_WIDTH-1:0]   mem_in_6_q1,
		output		[MEM_IN_6_DATA_WIDTH-1:0] 	mem_in_6_d1,
		
		output		[MEM_IN_7_ADDR_WIDTH-1:0] 	mem_in_7_addr1,
		output		 							mem_in_7_ce1,
		output		 							mem_in_7_we1,
		input 		[MEM_IN_7_DATA_WIDTH-1:0]   mem_in_7_q1,
		output		[MEM_IN_7_DATA_WIDTH-1:0] 	mem_in_7_d1,
		
		output		[MEM_IN_8_ADDR_WIDTH-1:0] 	mem_in_8_addr1,
		output		 							mem_in_8_ce1,
		output		 							mem_in_8_we1,
		input 		[MEM_IN_8_DATA_WIDTH-1:0]   mem_in_8_q1,
		output		[MEM_IN_8_DATA_WIDTH-1:0] 	mem_in_8_d1,
		
		output		[MEM_IN_9_ADDR_WIDTH-1:0] 	mem_in_9_addr1,
		output		 							mem_in_9_ce1,
		output		 							mem_in_9_we1,
		input 		[MEM_IN_9_DATA_WIDTH-1:0]   mem_in_9_q1,
		output		[MEM_IN_9_DATA_WIDTH-1:0] 	mem_in_9_d1,

		output		[MEM_IN_10_ADDR_WIDTH-1:0] 	mem_in_10_addr1,
		output		 							mem_in_10_ce1,
		output		 							mem_in_10_we1,
		input 		[MEM_IN_10_DATA_WIDTH-1:0]  mem_in_10_q1,
		output		[MEM_IN_10_DATA_WIDTH-1:0] 	mem_in_10_d1,

		output		[MEM_IN_11_ADDR_WIDTH-1:0] 	mem_in_11_addr1,
		output		 							mem_in_11_ce1,
		output		 							mem_in_11_we1,
		input 		[MEM_IN_11_DATA_WIDTH-1:0]  mem_in_11_q1,
		output		[MEM_IN_11_DATA_WIDTH-1:0] 	mem_in_11_d1,

		output		[MEM_IN_12_ADDR_WIDTH-1:0] 	mem_in_12_addr1,
		output		 							mem_in_12_ce1,
		output		 							mem_in_12_we1,
		input 		[MEM_IN_12_DATA_WIDTH-1:0]  mem_in_12_q1,
		output		[MEM_IN_12_DATA_WIDTH-1:0] 	mem_in_12_d1,

		output		[MEM_IN_13_ADDR_WIDTH-1:0] 	mem_in_13_addr1,
		output		 							mem_in_13_ce1,
		output		 							mem_in_13_we1,
		input 		[MEM_IN_13_DATA_WIDTH-1:0]  mem_in_13_q1,
		output		[MEM_IN_13_DATA_WIDTH-1:0] 	mem_in_13_d1,

		output		[MEM_IN_14_ADDR_WIDTH-1:0] 	mem_in_14_addr1,
		output		 							mem_in_14_ce1,
		output		 							mem_in_14_we1,
		input 		[MEM_IN_14_DATA_WIDTH-1:0]  mem_in_14_q1,
		output		[MEM_IN_14_DATA_WIDTH-1:0] 	mem_in_14_d1,

		output		[MEM_IN_15_ADDR_WIDTH-1:0] 	mem_in_15_addr1,
		output		 							mem_in_15_ce1,
		output		 							mem_in_15_we1,
		input 		[MEM_IN_15_DATA_WIDTH-1:0]  mem_in_15_q1,
		output		[MEM_IN_15_DATA_WIDTH-1:0] 	mem_in_15_d1,
		
		// Output Bram
		output		[MEM_OUT_0_ADDR_WIDTH-1:0] 	mem_out_0_addr1,
		output		 							mem_out_0_ce1,
		output		 							mem_out_0_we1,
		input 		[MEM_OUT_0_DATA_WIDTH-1:0]  mem_out_0_q1,
		output		[MEM_OUT_0_DATA_WIDTH-1:0] 	mem_out_0_d1,

		output		[MEM_OUT_1_ADDR_WIDTH-1:0] 	mem_out_1_addr1,
		output		 							mem_out_1_ce1,
		output		 							mem_out_1_we1,
		input 		[MEM_OUT_1_DATA_WIDTH-1:0]  mem_out_1_q1,
		output		[MEM_OUT_1_DATA_WIDTH-1:0] 	mem_out_1_d1,

		output		[MEM_OUT_2_ADDR_WIDTH-1:0] 	mem_out_2_addr1,
		output		 							mem_out_2_ce1,
		output		 							mem_out_2_we1,
		input 		[MEM_OUT_2_DATA_WIDTH-1:0]  mem_out_2_q1,
		output		[MEM_OUT_2_DATA_WIDTH-1:0] 	mem_out_2_d1,

		output		[MEM_OUT_3_ADDR_WIDTH-1:0] 	mem_out_3_addr1,
		output		 							mem_out_3_ce1,
		output		 							mem_out_3_we1,
		input 		[MEM_OUT_3_DATA_WIDTH-1:0]  mem_out_3_q1,
		output		[MEM_OUT_3_DATA_WIDTH-1:0] 	mem_out_3_d1,

		output		[MEM_OUT_4_ADDR_WIDTH-1:0] 	mem_out_4_addr1,
		output		 							mem_out_4_ce1,
		output		 							mem_out_4_we1,
		input 		[MEM_OUT_4_DATA_WIDTH-1:0]  mem_out_4_q1,
		output		[MEM_OUT_4_DATA_WIDTH-1:0] 	mem_out_4_d1,

		output		[MEM_OUT_5_ADDR_WIDTH-1:0] 	mem_out_5_addr1,
		output		 							mem_out_5_ce1,
		output		 							mem_out_5_we1,
		input 		[MEM_OUT_5_DATA_WIDTH-1:0]  mem_out_5_q1,
		output		[MEM_OUT_5_DATA_WIDTH-1:0] 	mem_out_5_d1,

		output		[MEM_OUT_6_ADDR_WIDTH-1:0] 	mem_out_6_addr1,
		output		 							mem_out_6_ce1,
		output		 							mem_out_6_we1,
		input 		[MEM_OUT_6_DATA_WIDTH-1:0]  mem_out_6_q1,
		output		[MEM_OUT_6_DATA_WIDTH-1:0] 	mem_out_6_d1,

		output		[MEM_OUT_7_ADDR_WIDTH-1:0] 	mem_out_7_addr1,
		output		 							mem_out_7_ce1,
		output		 							mem_out_7_we1,
		input 		[MEM_OUT_7_DATA_WIDTH-1:0]  mem_out_7_q1,
		output		[MEM_OUT_7_DATA_WIDTH-1:0] 	mem_out_7_d1,

		output		[MEM_OUT_8_ADDR_WIDTH-1:0] 	mem_out_8_addr1,
		output		 							mem_out_8_ce1,
		output		 							mem_out_8_we1,
		input 		[MEM_OUT_8_DATA_WIDTH-1:0]  mem_out_8_q1,
		output		[MEM_OUT_8_DATA_WIDTH-1:0] 	mem_out_8_d1,

		output		[MEM_OUT_9_ADDR_WIDTH-1:0] 	mem_out_9_addr1,
		output		 							mem_out_9_ce1,
		output		 							mem_out_9_we1,
		input 		[MEM_OUT_9_DATA_WIDTH-1:0]  mem_out_9_q1,
		output		[MEM_OUT_9_DATA_WIDTH-1:0] 	mem_out_9_d1,

		output		[MEM_OUT_10_ADDR_WIDTH-1:0] mem_out_10_addr1,
		output		 							mem_out_10_ce1,
		output		 							mem_out_10_we1,
		input 		[MEM_OUT_10_DATA_WIDTH-1:0] mem_out_10_q1,
		output		[MEM_OUT_10_DATA_WIDTH-1:0] mem_out_10_d1,

		output		[MEM_OUT_11_ADDR_WIDTH-1:0] mem_out_11_addr1,
		output		 							mem_out_11_ce1,
		output		 							mem_out_11_we1,
		input 		[MEM_OUT_11_DATA_WIDTH-1:0] mem_out_11_q1,
		output		[MEM_OUT_11_DATA_WIDTH-1:0] mem_out_11_d1,

		output		[MEM_OUT_12_ADDR_WIDTH-1:0] mem_out_12_addr1,
		output		 							mem_out_12_ce1,
		output		 							mem_out_12_we1,
		input 		[MEM_OUT_12_DATA_WIDTH-1:0] mem_out_12_q1,
		output		[MEM_OUT_12_DATA_WIDTH-1:0] mem_out_12_d1,

		output		[MEM_OUT_13_ADDR_WIDTH-1:0] mem_out_13_addr1,
		output		 							mem_out_13_ce1,
		output		 							mem_out_13_we1,
		input 		[MEM_OUT_13_DATA_WIDTH-1:0] mem_out_13_q1,
		output		[MEM_OUT_13_DATA_WIDTH-1:0] mem_out_13_d1,

		output		[MEM_OUT_14_ADDR_WIDTH-1:0] mem_out_14_addr1,
		output		 							mem_out_14_ce1,
		output		 							mem_out_14_we1,
		input 		[MEM_OUT_14_DATA_WIDTH-1:0] mem_out_14_q1,
		output		[MEM_OUT_14_DATA_WIDTH-1:0] mem_out_14_d1,

		output		[MEM_OUT_15_ADDR_WIDTH-1:0] mem_out_15_addr1,
		output		 							mem_out_15_ce1,
		output		 							mem_out_15_we1,
		input 		[MEM_OUT_15_DATA_WIDTH-1:0] mem_out_15_q1,
		output		[MEM_OUT_15_DATA_WIDTH-1:0] mem_out_15_d1,

		output		[MEM_OUT_16_ADDR_WIDTH-1:0] mem_out_16_addr1,
		output		 							mem_out_16_ce1,
		output		 							mem_out_16_we1,
		input 		[MEM_OUT_16_DATA_WIDTH-1:0] mem_out_16_q1,
		output		[MEM_OUT_16_DATA_WIDTH-1:0] mem_out_16_d1,

		output		[MEM_OUT_17_ADDR_WIDTH-1:0] mem_out_17_addr1,
		output		 							mem_out_17_ce1,
		output		 							mem_out_17_we1,
		input 		[MEM_OUT_17_DATA_WIDTH-1:0] mem_out_17_q1,
		output		[MEM_OUT_17_DATA_WIDTH-1:0] mem_out_17_d1,

		input		[C_S00_AXI_DATA_WIDTH-1:0]	fsm_status_reg_in,
		output		[C_S00_AXI_DATA_WIDTH-1:0]	fsm_status_reg_out,


		// User ports ends
		// Do not modify the ports beyond this line


		// Ports of Axi Slave Bus Interface S00_AXI
		input wire  s00_axi_aclk,
		input wire  s00_axi_aresetn,
		input wire [C_S00_AXI_ADDR_WIDTH-1 : 0] s00_axi_awaddr,
		input wire [2 : 0] s00_axi_awprot,
		input wire  s00_axi_awvalid,
		output wire  s00_axi_awready,
		input wire [C_S00_AXI_DATA_WIDTH-1 : 0] s00_axi_wdata,
		input wire [(C_S00_AXI_DATA_WIDTH/8)-1 : 0] s00_axi_wstrb,
		input wire  s00_axi_wvalid,
		output wire  s00_axi_wready,
		output wire [1 : 0] s00_axi_bresp,
		output wire  s00_axi_bvalid,
		input wire  s00_axi_bready,
		input wire [C_S00_AXI_ADDR_WIDTH-1 : 0] s00_axi_araddr,
		input wire [2 : 0] s00_axi_arprot,
		input wire  s00_axi_arvalid,
		output wire  s00_axi_arready,
		output wire [C_S00_AXI_DATA_WIDTH-1 : 0] s00_axi_rdata,
		output wire [1 : 0] s00_axi_rresp,
		output wire  s00_axi_rvalid,
		input wire  s00_axi_rready
	);

	// Instantiation of Axi Bus Interface S00_AXI
	myip_v1_0_S00_AXI # (
		.CNT_BIT(CNT_BIT),
		
		.MEM_IN_0_DATA_WIDTH(MEM_IN_0_DATA_WIDTH),
		.MEM_IN_0_ADDR_WIDTH(MEM_IN_0_ADDR_WIDTH),
		.MEM_IN_1_DATA_WIDTH(MEM_IN_1_DATA_WIDTH),
		.MEM_IN_1_ADDR_WIDTH(MEM_IN_1_ADDR_WIDTH),
		.MEM_IN_2_DATA_WIDTH(MEM_IN_2_DATA_WIDTH),
		.MEM_IN_2_ADDR_WIDTH(MEM_IN_2_ADDR_WIDTH),
		.MEM_IN_3_DATA_WIDTH(MEM_IN_3_DATA_WIDTH),
		.MEM_IN_3_ADDR_WIDTH(MEM_IN_3_ADDR_WIDTH),
		.MEM_IN_4_DATA_WIDTH(MEM_IN_4_DATA_WIDTH),
		.MEM_IN_4_ADDR_WIDTH(MEM_IN_4_ADDR_WIDTH),
		.MEM_IN_5_DATA_WIDTH(MEM_IN_5_DATA_WIDTH),
		.MEM_IN_5_ADDR_WIDTH(MEM_IN_5_ADDR_WIDTH),
		.MEM_IN_6_DATA_WIDTH(MEM_IN_6_DATA_WIDTH),
		.MEM_IN_6_ADDR_WIDTH(MEM_IN_6_ADDR_WIDTH),
		.MEM_IN_7_DATA_WIDTH(MEM_IN_7_DATA_WIDTH),
		.MEM_IN_7_ADDR_WIDTH(MEM_IN_7_ADDR_WIDTH),
		.MEM_IN_8_DATA_WIDTH(MEM_IN_8_DATA_WIDTH),
		.MEM_IN_8_ADDR_WIDTH(MEM_IN_8_ADDR_WIDTH),
		.MEM_IN_9_DATA_WIDTH(MEM_IN_9_DATA_WIDTH),
		.MEM_IN_9_ADDR_WIDTH(MEM_IN_9_ADDR_WIDTH),
		.MEM_IN_10_DATA_WIDTH(MEM_IN_10_DATA_WIDTH),
		.MEM_IN_10_ADDR_WIDTH(MEM_IN_10_ADDR_WIDTH),
		.MEM_IN_11_DATA_WIDTH(MEM_IN_11_DATA_WIDTH),
		.MEM_IN_11_ADDR_WIDTH(MEM_IN_11_ADDR_WIDTH),
		.MEM_IN_12_DATA_WIDTH(MEM_IN_12_DATA_WIDTH),
		.MEM_IN_12_ADDR_WIDTH(MEM_IN_12_ADDR_WIDTH),
		.MEM_IN_13_DATA_WIDTH(MEM_IN_13_DATA_WIDTH),
		.MEM_IN_13_ADDR_WIDTH(MEM_IN_13_ADDR_WIDTH),
		.MEM_IN_14_DATA_WIDTH(MEM_IN_14_DATA_WIDTH),
		.MEM_IN_14_ADDR_WIDTH(MEM_IN_14_ADDR_WIDTH),
		.MEM_IN_15_DATA_WIDTH(MEM_IN_15_DATA_WIDTH),
		.MEM_IN_15_ADDR_WIDTH(MEM_IN_15_ADDR_WIDTH),

		.MEM_OUT_0_DATA_WIDTH(MEM_OUT_0_DATA_WIDTH),
		.MEM_OUT_0_ADDR_WIDTH(MEM_OUT_0_ADDR_WIDTH),
		.MEM_OUT_1_DATA_WIDTH(MEM_OUT_1_DATA_WIDTH),
		.MEM_OUT_1_ADDR_WIDTH(MEM_OUT_1_ADDR_WIDTH),
		.MEM_OUT_2_DATA_WIDTH(MEM_OUT_2_DATA_WIDTH),
		.MEM_OUT_2_ADDR_WIDTH(MEM_OUT_2_ADDR_WIDTH),
		.MEM_OUT_3_DATA_WIDTH(MEM_OUT_3_DATA_WIDTH),
		.MEM_OUT_3_ADDR_WIDTH(MEM_OUT_3_ADDR_WIDTH),
		.MEM_OUT_4_DATA_WIDTH(MEM_OUT_4_DATA_WIDTH),
		.MEM_OUT_4_ADDR_WIDTH(MEM_OUT_4_ADDR_WIDTH),
		.MEM_OUT_5_DATA_WIDTH(MEM_OUT_5_DATA_WIDTH),
		.MEM_OUT_5_ADDR_WIDTH(MEM_OUT_5_ADDR_WIDTH),
		.MEM_OUT_6_DATA_WIDTH(MEM_OUT_6_DATA_WIDTH),
		.MEM_OUT_6_ADDR_WIDTH(MEM_OUT_6_ADDR_WIDTH),
		.MEM_OUT_7_DATA_WIDTH(MEM_OUT_7_DATA_WIDTH),
		.MEM_OUT_7_ADDR_WIDTH(MEM_OUT_7_ADDR_WIDTH),
		.MEM_OUT_8_DATA_WIDTH(MEM_OUT_8_DATA_WIDTH),
		.MEM_OUT_8_ADDR_WIDTH(MEM_OUT_8_ADDR_WIDTH),
		.MEM_OUT_9_DATA_WIDTH(MEM_OUT_9_DATA_WIDTH),
		.MEM_OUT_9_ADDR_WIDTH(MEM_OUT_9_ADDR_WIDTH),
		.MEM_OUT_10_DATA_WIDTH(MEM_OUT_10_DATA_WIDTH),
		.MEM_OUT_10_ADDR_WIDTH(MEM_OUT_10_ADDR_WIDTH),
		.MEM_OUT_11_DATA_WIDTH(MEM_OUT_11_DATA_WIDTH),
		.MEM_OUT_11_ADDR_WIDTH(MEM_OUT_11_ADDR_WIDTH),
		.MEM_OUT_12_DATA_WIDTH(MEM_OUT_12_DATA_WIDTH),
		.MEM_OUT_12_ADDR_WIDTH(MEM_OUT_12_ADDR_WIDTH),
		.MEM_OUT_13_DATA_WIDTH(MEM_OUT_13_DATA_WIDTH),
		.MEM_OUT_13_ADDR_WIDTH(MEM_OUT_13_ADDR_WIDTH),
		.MEM_OUT_14_DATA_WIDTH(MEM_OUT_14_DATA_WIDTH),
		.MEM_OUT_14_ADDR_WIDTH(MEM_OUT_14_ADDR_WIDTH),
		.MEM_OUT_15_DATA_WIDTH(MEM_OUT_15_DATA_WIDTH),
		.MEM_OUT_15_ADDR_WIDTH(MEM_OUT_15_ADDR_WIDTH),
		.MEM_OUT_16_DATA_WIDTH(MEM_OUT_16_DATA_WIDTH),
		.MEM_OUT_16_ADDR_WIDTH(MEM_OUT_16_ADDR_WIDTH),
		.MEM_OUT_17_DATA_WIDTH(MEM_OUT_17_DATA_WIDTH),
		.MEM_OUT_17_ADDR_WIDTH(MEM_OUT_17_ADDR_WIDTH),

		.C_S_AXI_DATA_WIDTH(C_S00_AXI_DATA_WIDTH),
		.C_S_AXI_ADDR_WIDTH(C_S00_AXI_ADDR_WIDTH)
	) myip_v1_0_S00_AXI_inst (
		.mem_in_0_addr1(mem_in_0_addr1),
		.mem_in_0_ce1(mem_in_0_ce1),
		.mem_in_0_we1(mem_in_0_we1),
		.mem_in_0_q1(mem_in_0_q1),
		.mem_in_0_d1(mem_in_0_d1),
		.mem_in_1_addr1(mem_in_1_addr1),
		.mem_in_1_ce1(mem_in_1_ce1),
		.mem_in_1_we1(mem_in_1_we1),
		.mem_in_1_q1(mem_in_1_q1),
		.mem_in_1_d1(mem_in_1_d1),
		.mem_in_2_addr1(mem_in_2_addr1),
		.mem_in_2_ce1(mem_in_2_ce1),
		.mem_in_2_we1(mem_in_2_we1),
		.mem_in_2_q1(mem_in_2_q1),
		.mem_in_2_d1(mem_in_2_d1),
		.mem_in_3_addr1(mem_in_3_addr1),
		.mem_in_3_ce1(mem_in_3_ce1),
		.mem_in_3_we1(mem_in_3_we1),
		.mem_in_3_q1(mem_in_3_q1),
		.mem_in_3_d1(mem_in_3_d1),
		.mem_in_4_addr1(mem_in_4_addr1),
		.mem_in_4_ce1(mem_in_4_ce1),
		.mem_in_4_we1(mem_in_4_we1),
		.mem_in_4_q1(mem_in_4_q1),
		.mem_in_4_d1(mem_in_4_d1),
		.mem_in_5_addr1(mem_in_5_addr1),
		.mem_in_5_ce1(mem_in_5_ce1),
		.mem_in_5_we1(mem_in_5_we1),
		.mem_in_5_q1(mem_in_5_q1),
		.mem_in_5_d1(mem_in_5_d1),
		.mem_in_6_addr1(mem_in_6_addr1),
		.mem_in_6_ce1(mem_in_6_ce1),
		.mem_in_6_we1(mem_in_6_we1),
		.mem_in_6_q1(mem_in_6_q1),
		.mem_in_6_d1(mem_in_6_d1),
		.mem_in_7_addr1(mem_in_7_addr1),
		.mem_in_7_ce1(mem_in_7_ce1),
		.mem_in_7_we1(mem_in_7_we1),
		.mem_in_7_q1(mem_in_7_q1),
		.mem_in_7_d1(mem_in_7_d1),
		.mem_in_8_addr1(mem_in_8_addr1),
		.mem_in_8_ce1(mem_in_8_ce1),
		.mem_in_8_we1(mem_in_8_we1),
		.mem_in_8_q1(mem_in_8_q1),
		.mem_in_8_d1(mem_in_8_d1),
		.mem_in_9_addr1(mem_in_9_addr1),
		.mem_in_9_ce1(mem_in_9_ce1),
		.mem_in_9_we1(mem_in_9_we1),
		.mem_in_9_q1(mem_in_9_q1),
		.mem_in_9_d1(mem_in_9_d1),
		.mem_in_10_addr1(mem_in_10_addr1),
		.mem_in_10_ce1(mem_in_10_ce1),
		.mem_in_10_we1(mem_in_10_we1),
		.mem_in_10_q1(mem_in_10_q1),
		.mem_in_10_d1(mem_in_10_d1),
		.mem_in_11_addr1(mem_in_11_addr1),
		.mem_in_11_ce1(mem_in_11_ce1),
		.mem_in_11_we1(mem_in_11_we1),
		.mem_in_11_q1(mem_in_11_q1),
		.mem_in_11_d1(mem_in_11_d1),
		.mem_in_12_addr1(mem_in_12_addr1),
		.mem_in_12_ce1(mem_in_12_ce1),
		.mem_in_12_we1(mem_in_12_we1),
		.mem_in_12_q1(mem_in_12_q1),
		.mem_in_12_d1(mem_in_12_d1),
		.mem_in_13_addr1(mem_in_13_addr1),
		.mem_in_13_ce1(mem_in_13_ce1),
		.mem_in_13_we1(mem_in_13_we1),
		.mem_in_13_q1(mem_in_13_q1),
		.mem_in_13_d1(mem_in_13_d1),
		.mem_in_14_addr1(mem_in_14_addr1),
		.mem_in_14_ce1(mem_in_14_ce1),
		.mem_in_14_we1(mem_in_14_we1),
		.mem_in_14_q1(mem_in_14_q1),
		.mem_in_14_d1(mem_in_14_d1),
		.mem_in_15_addr1(mem_in_15_addr1),
		.mem_in_15_ce1(mem_in_15_ce1),
		.mem_in_15_we1(mem_in_15_we1),
		.mem_in_15_q1(mem_in_15_q1),
		.mem_in_15_d1(mem_in_15_d1),

		.mem_out_0_addr1(mem_out_0_addr1),
		.mem_out_0_ce1(mem_out_0_ce1),
		.mem_out_0_we1(mem_out_0_we1),
		.mem_out_0_q1(mem_out_0_q1),
		.mem_out_0_d1(mem_out_0_d1),
		.mem_out_1_addr1(mem_out_1_addr1),
		.mem_out_1_ce1(mem_out_1_ce1),
		.mem_out_1_we1(mem_out_1_we1),
		.mem_out_1_q1(mem_out_1_q1),
		.mem_out_1_d1(mem_out_1_d1),
		.mem_out_2_addr1(mem_out_2_addr1),
		.mem_out_2_ce1(mem_out_2_ce1),
		.mem_out_2_we1(mem_out_2_we1),
		.mem_out_2_q1(mem_out_2_q1),
		.mem_out_2_d1(mem_out_2_d1),
		.mem_out_3_addr1(mem_out_3_addr1),
		.mem_out_3_ce1(mem_out_3_ce1),
		.mem_out_3_we1(mem_out_3_we1),
		.mem_out_3_q1(mem_out_3_q1),
		.mem_out_3_d1(mem_out_3_d1),
		.mem_out_4_addr1(mem_out_4_addr1),
		.mem_out_4_ce1(mem_out_4_ce1),
		.mem_out_4_we1(mem_out_4_we1),
		.mem_out_4_q1(mem_out_4_q1),
		.mem_out_4_d1(mem_out_4_d1),
		.mem_out_5_addr1(mem_out_5_addr1),
		.mem_out_5_ce1(mem_out_5_ce1),
		.mem_out_5_we1(mem_out_5_we1),
		.mem_out_5_q1(mem_out_5_q1),
		.mem_out_5_d1(mem_out_5_d1),
		.mem_out_6_addr1(mem_out_6_addr1),
		.mem_out_6_ce1(mem_out_6_ce1),
		.mem_out_6_we1(mem_out_6_we1),
		.mem_out_6_q1(mem_out_6_q1),
		.mem_out_6_d1(mem_out_6_d1),
		.mem_out_7_addr1(mem_out_7_addr1),
		.mem_out_7_ce1(mem_out_7_ce1),
		.mem_out_7_we1(mem_out_7_we1),
		.mem_out_7_q1(mem_out_7_q1),
		.mem_out_7_d1(mem_out_7_d1),
		.mem_out_8_addr1(mem_out_8_addr1),
		.mem_out_8_ce1(mem_out_8_ce1),
		.mem_out_8_we1(mem_out_8_we1),
		.mem_out_8_q1(mem_out_8_q1),
		.mem_out_8_d1(mem_out_8_d1),
		.mem_out_9_addr1(mem_out_9_addr1),
		.mem_out_9_ce1(mem_out_9_ce1),
		.mem_out_9_we1(mem_out_9_we1),
		.mem_out_9_q1(mem_out_9_q1),
		.mem_out_9_d1(mem_out_9_d1),
		.mem_out_10_addr1(mem_out_10_addr1),
		.mem_out_10_ce1(mem_out_10_ce1),
		.mem_out_10_we1(mem_out_10_we1),
		.mem_out_10_q1(mem_out_10_q1),
		.mem_out_10_d1(mem_out_10_d1),
		.mem_out_11_addr1(mem_out_11_addr1),
		.mem_out_11_ce1(mem_out_11_ce1),
		.mem_out_11_we1(mem_out_11_we1),
		.mem_out_11_q1(mem_out_11_q1),
		.mem_out_11_d1(mem_out_11_d1),
		.mem_out_12_addr1(mem_out_12_addr1),
		.mem_out_12_ce1(mem_out_12_ce1),
		.mem_out_12_we1(mem_out_12_we1),
		.mem_out_12_q1(mem_out_12_q1),
		.mem_out_12_d1(mem_out_12_d1),
		.mem_out_13_addr1(mem_out_13_addr1),
		.mem_out_13_ce1(mem_out_13_ce1),
		.mem_out_13_we1(mem_out_13_we1),
		.mem_out_13_q1(mem_out_13_q1),
		.mem_out_13_d1(mem_out_13_d1),
		.mem_out_14_addr1(mem_out_14_addr1),
		.mem_out_14_ce1(mem_out_14_ce1),
		.mem_out_14_we1(mem_out_14_we1),
		.mem_out_14_q1(mem_out_14_q1),
		.mem_out_14_d1(mem_out_14_d1),
		.mem_out_15_addr1(mem_out_15_addr1),
		.mem_out_15_ce1(mem_out_15_ce1),
		.mem_out_15_we1(mem_out_15_we1),
		.mem_out_15_q1(mem_out_15_q1),
		.mem_out_15_d1(mem_out_15_d1),
		.mem_out_16_addr1(mem_out_16_addr1),
		.mem_out_16_ce1(mem_out_16_ce1),
		.mem_out_16_we1(mem_out_16_we1),
		.mem_out_16_q1(mem_out_16_q1),
		.mem_out_16_d1(mem_out_16_d1),
		.mem_out_17_addr1(mem_out_17_addr1),
		.mem_out_17_ce1(mem_out_17_ce1),
		.mem_out_17_we1(mem_out_17_we1),
		.mem_out_17_q1(mem_out_17_q1),
		.mem_out_17_d1(mem_out_17_d1),
		.fsm_status_reg_in(fsm_status_reg_in),
		.fsm_status_reg_out(fsm_status_reg_out),

		.S_AXI_ACLK(s00_axi_aclk),
		.S_AXI_ARESETN(s00_axi_aresetn),
		.S_AXI_AWADDR(s00_axi_awaddr),
		.S_AXI_AWPROT(s00_axi_awprot),
		.S_AXI_AWVALID(s00_axi_awvalid),
		.S_AXI_AWREADY(s00_axi_awready),
		.S_AXI_WDATA(s00_axi_wdata),
		.S_AXI_WSTRB(s00_axi_wstrb),
		.S_AXI_WVALID(s00_axi_wvalid),
		.S_AXI_WREADY(s00_axi_wready),
		.S_AXI_BRESP(s00_axi_bresp),
		.S_AXI_BVALID(s00_axi_bvalid),
		.S_AXI_BREADY(s00_axi_bready),
		.S_AXI_ARADDR(s00_axi_araddr),
		.S_AXI_ARPROT(s00_axi_arprot),
		.S_AXI_ARVALID(s00_axi_arvalid),
		.S_AXI_ARREADY(s00_axi_arready),
		.S_AXI_RDATA(s00_axi_rdata),
		.S_AXI_RRESP(s00_axi_rresp),
		.S_AXI_RVALID(s00_axi_rvalid),
		.S_AXI_RREADY(s00_axi_rready)
	);

	// Add user logic here

	// User logic ends

	endmodule
